// mysystem.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module mysystem (
		input  wire        alt_vip_itc_0_clocked_video_vid_clk,       //  alt_vip_itc_0_clocked_video.vid_clk
		output wire [31:0] alt_vip_itc_0_clocked_video_vid_data,      //                             .vid_data
		output wire        alt_vip_itc_0_clocked_video_underflow,     //                             .underflow
		output wire        alt_vip_itc_0_clocked_video_vid_datavalid, //                             .vid_datavalid
		output wire        alt_vip_itc_0_clocked_video_vid_v_sync,    //                             .vid_v_sync
		output wire        alt_vip_itc_0_clocked_video_vid_h_sync,    //                             .vid_h_sync
		output wire        alt_vip_itc_0_clocked_video_vid_f,         //                             .vid_f
		output wire        alt_vip_itc_0_clocked_video_vid_h,         //                             .vid_h
		output wire        alt_vip_itc_0_clocked_video_vid_v,         //                             .vid_v
		output wire        clk_65_clk,                                //                       clk_65.clk
		input  wire        donesig_export,                            //                      donesig.export
		output wire        hps_0_h2f_reset_reset_n,                   //              hps_0_h2f_reset.reset_n
		inout  wire        hps_io_hps_io_sdio_inst_CMD,               //                       hps_io.hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,                //                             .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,                //                             .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,               //                             .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,                //                             .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,                //                             .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,                //                             .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,                //                             .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,                //                             .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,                //                             .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,                //                             .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,                //                             .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,                //                             .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,                //                             .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,               //                             .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,               //                             .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,               //                             .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,               //                             .hps_io_usb1_inst_NXT
		input  wire        hps_io_hps_io_uart0_inst_RX,               //                             .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,               //                             .hps_io_uart0_inst_TX
		output wire [9:0]  led_external_connection_export,            //      led_external_connection.export
		output wire [14:0] memory_mem_a,                              //                       memory.mem_a
		output wire [2:0]  memory_mem_ba,                             //                             .mem_ba
		output wire        memory_mem_ck,                             //                             .mem_ck
		output wire        memory_mem_ck_n,                           //                             .mem_ck_n
		output wire        memory_mem_cke,                            //                             .mem_cke
		output wire        memory_mem_cs_n,                           //                             .mem_cs_n
		output wire        memory_mem_ras_n,                          //                             .mem_ras_n
		output wire        memory_mem_cas_n,                          //                             .mem_cas_n
		output wire        memory_mem_we_n,                           //                             .mem_we_n
		output wire        memory_mem_reset_n,                        //                             .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                             //                             .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                            //                             .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                          //                             .mem_dqs_n
		output wire        memory_mem_odt,                            //                             .mem_odt
		output wire [3:0]  memory_mem_dm,                             //                             .mem_dm
		input  wire        memory_oct_rzqin,                          //                             .oct_rzqin
		output wire        sdram_clk_clk,                             //                    sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                           //                   sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                             //                             .ba
		output wire        sdram_wire_cas_n,                          //                             .cas_n
		output wire        sdram_wire_cke,                            //                             .cke
		output wire        sdram_wire_cs_n,                           //                             .cs_n
		inout  wire [15:0] sdram_wire_dq,                             //                             .dq
		output wire [1:0]  sdram_wire_dqm,                            //                             .dqm
		output wire        sdram_wire_ras_n,                          //                             .ras_n
		output wire        sdram_wire_we_n,                           //                             .we_n
		output wire [3:0]  sdramstartstop_readdata,                   //               sdramstartstop.readdata
		input  wire        sdramstartstop_beginbursttransfer,         //                             .beginbursttransfer
		output wire        sdramstartstop_writeresponsevalid_n,       //                             .writeresponsevalid_n
		output wire        startsig_export,                           //                     startsig.export
		input  wire [9:0]  switches_external_connection_export,       // switches_external_connection.export
		input  wire        system_ref_clk_clk,                        //               system_ref_clk.clk
		input  wire        system_ref_reset_reset                     //             system_ref_reset.reset
	);

	wire          alt_vip_vfr_0_avalon_streaming_source_valid;                 // alt_vip_vfr_0:dout_valid -> alt_vip_itc_0:is_valid
	wire   [31:0] alt_vip_vfr_0_avalon_streaming_source_data;                  // alt_vip_vfr_0:dout_data -> alt_vip_itc_0:is_data
	wire          alt_vip_vfr_0_avalon_streaming_source_ready;                 // alt_vip_itc_0:is_ready -> alt_vip_vfr_0:dout_ready
	wire          alt_vip_vfr_0_avalon_streaming_source_startofpacket;         // alt_vip_vfr_0:dout_startofpacket -> alt_vip_itc_0:is_sop
	wire          alt_vip_vfr_0_avalon_streaming_source_endofpacket;           // alt_vip_vfr_0:dout_endofpacket -> alt_vip_itc_0:is_eop
	wire          pll_0_outclk0_clk;                                           // pll_0:outclk_0 -> [alt_vip_itc_0:is_clk, alt_vip_vfr_0:clock, mm_interconnect_2:pll_0_outclk0_clk, rst_controller:clk]
	wire          sys_clk_sys_clk_clk;                                         // sys_clk:sys_clk_clk -> [alt_vip_vfr_0:master_clock, doneSignal:clk, hps_0:f2h_axi_clk, hps_0:h2f_axi_clk, hps_0:h2f_lw_axi_clk, jtag_uart_0:clk, led:clk, mm_interconnect_0:sys_clk_sys_clk_clk, mm_interconnect_1:sys_clk_sys_clk_clk, mm_interconnect_2:sys_clk_sys_clk_clk, pll_0:refclk, pll_1:refclk, rst_controller_001:clk, rst_controller_002:clk, sdram_controller:clk, sdram_master_0:clk, startSignal:clk, switches:clk, sysid_qsys_0:clock]
	wire          sys_clk_reset_source_reset;                                  // sys_clk:reset_source_reset -> [pll_0:rst, pll_1:rst, rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire  [127:0] alt_vip_vfr_0_avalon_master_readdata;                        // mm_interconnect_0:alt_vip_vfr_0_avalon_master_readdata -> alt_vip_vfr_0:master_readdata
	wire          alt_vip_vfr_0_avalon_master_waitrequest;                     // mm_interconnect_0:alt_vip_vfr_0_avalon_master_waitrequest -> alt_vip_vfr_0:master_waitrequest
	wire   [31:0] alt_vip_vfr_0_avalon_master_address;                         // alt_vip_vfr_0:master_address -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_address
	wire          alt_vip_vfr_0_avalon_master_read;                            // alt_vip_vfr_0:master_read -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_read
	wire          alt_vip_vfr_0_avalon_master_readdatavalid;                   // mm_interconnect_0:alt_vip_vfr_0_avalon_master_readdatavalid -> alt_vip_vfr_0:master_readdatavalid
	wire    [5:0] alt_vip_vfr_0_avalon_master_burstcount;                      // alt_vip_vfr_0:master_burstcount -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_burstcount
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_awburst;               // mm_interconnect_0:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire    [4:0] mm_interconnect_0_hps_0_f2h_axi_slave_awuser;                // mm_interconnect_0:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_arlen;                 // mm_interconnect_0:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire   [15:0] mm_interconnect_0_hps_0_f2h_axi_slave_wstrb;                 // mm_interconnect_0:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_wready;                // hps_0:f2h_WREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_wready
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_rid;                   // hps_0:f2h_RID -> mm_interconnect_0:hps_0_f2h_axi_slave_rid
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_rready;                // mm_interconnect_0:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_awlen;                 // mm_interconnect_0:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_wid;                   // mm_interconnect_0:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_arcache;               // mm_interconnect_0:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_wvalid;                // mm_interconnect_0:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire   [31:0] mm_interconnect_0_hps_0_f2h_axi_slave_araddr;                // mm_interconnect_0:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_arprot;                // mm_interconnect_0:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_awprot;                // mm_interconnect_0:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire  [127:0] mm_interconnect_0_hps_0_f2h_axi_slave_wdata;                 // mm_interconnect_0:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_arvalid;               // mm_interconnect_0:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_awcache;               // mm_interconnect_0:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_arid;                  // mm_interconnect_0:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_arlock;                // mm_interconnect_0:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_awlock;                // mm_interconnect_0:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire   [31:0] mm_interconnect_0_hps_0_f2h_axi_slave_awaddr;                // mm_interconnect_0:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_bresp;                 // hps_0:f2h_BRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_bresp
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_arready;               // hps_0:f2h_ARREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_arready
	wire  [127:0] mm_interconnect_0_hps_0_f2h_axi_slave_rdata;                 // hps_0:f2h_RDATA -> mm_interconnect_0:hps_0_f2h_axi_slave_rdata
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_awready;               // hps_0:f2h_AWREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_awready
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_arburst;               // mm_interconnect_0:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_arsize;                // mm_interconnect_0:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_bready;                // mm_interconnect_0:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_rlast;                 // hps_0:f2h_RLAST -> mm_interconnect_0:hps_0_f2h_axi_slave_rlast
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_wlast;                 // mm_interconnect_0:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_rresp;                 // hps_0:f2h_RRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_rresp
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_awid;                  // mm_interconnect_0:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_bid;                   // hps_0:f2h_BID -> mm_interconnect_0:hps_0_f2h_axi_slave_bid
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_bvalid;                // hps_0:f2h_BVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_bvalid
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_awsize;                // mm_interconnect_0:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_awvalid;               // mm_interconnect_0:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire    [4:0] mm_interconnect_0_hps_0_f2h_axi_slave_aruser;                // mm_interconnect_0:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_rvalid;                // hps_0:f2h_RVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_rvalid
	wire          sdram_master_0_avalon_master_chipselect;                     // sdram_master_0:chipselect -> mm_interconnect_1:sdram_master_0_avalon_master_chipselect
	wire          sdram_master_0_avalon_master_waitrequest;                    // mm_interconnect_1:sdram_master_0_avalon_master_waitrequest -> sdram_master_0:waitrequest
	wire   [15:0] sdram_master_0_avalon_master_readdata;                       // mm_interconnect_1:sdram_master_0_avalon_master_readdata -> sdram_master_0:readdata
	wire          sdram_master_0_avalon_master_read;                           // sdram_master_0:read_n -> mm_interconnect_1:sdram_master_0_avalon_master_read
	wire   [31:0] sdram_master_0_avalon_master_address;                        // sdram_master_0:address -> mm_interconnect_1:sdram_master_0_avalon_master_address
	wire    [1:0] sdram_master_0_avalon_master_byteenable;                     // sdram_master_0:byteenable -> mm_interconnect_1:sdram_master_0_avalon_master_byteenable
	wire          sdram_master_0_avalon_master_readdatavalid;                  // mm_interconnect_1:sdram_master_0_avalon_master_readdatavalid -> sdram_master_0:readdatavalid
	wire          sdram_master_0_avalon_master_write;                          // sdram_master_0:write_n -> mm_interconnect_1:sdram_master_0_avalon_master_write
	wire   [15:0] sdram_master_0_avalon_master_writedata;                      // sdram_master_0:writedata -> mm_interconnect_1:sdram_master_0_avalon_master_writedata
	wire    [1:0] hps_0_h2f_axi_master_awburst;                                // hps_0:h2f_AWBURST -> mm_interconnect_1:hps_0_h2f_axi_master_awburst
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                  // hps_0:h2f_ARLEN -> mm_interconnect_1:hps_0_h2f_axi_master_arlen
	wire    [7:0] hps_0_h2f_axi_master_wstrb;                                  // hps_0:h2f_WSTRB -> mm_interconnect_1:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_wready;                                 // mm_interconnect_1:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [11:0] hps_0_h2f_axi_master_rid;                                    // mm_interconnect_1:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_rready;                                 // hps_0:h2f_RREADY -> mm_interconnect_1:hps_0_h2f_axi_master_rready
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                  // hps_0:h2f_AWLEN -> mm_interconnect_1:hps_0_h2f_axi_master_awlen
	wire   [11:0] hps_0_h2f_axi_master_wid;                                    // hps_0:h2f_WID -> mm_interconnect_1:hps_0_h2f_axi_master_wid
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                // hps_0:h2f_ARCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_arcache
	wire          hps_0_h2f_axi_master_wvalid;                                 // hps_0:h2f_WVALID -> mm_interconnect_1:hps_0_h2f_axi_master_wvalid
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                 // hps_0:h2f_ARADDR -> mm_interconnect_1:hps_0_h2f_axi_master_araddr
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                 // hps_0:h2f_ARPROT -> mm_interconnect_1:hps_0_h2f_axi_master_arprot
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                 // hps_0:h2f_AWPROT -> mm_interconnect_1:hps_0_h2f_axi_master_awprot
	wire   [63:0] hps_0_h2f_axi_master_wdata;                                  // hps_0:h2f_WDATA -> mm_interconnect_1:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_arvalid;                                // hps_0:h2f_ARVALID -> mm_interconnect_1:hps_0_h2f_axi_master_arvalid
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                // hps_0:h2f_AWCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_awcache
	wire   [11:0] hps_0_h2f_axi_master_arid;                                   // hps_0:h2f_ARID -> mm_interconnect_1:hps_0_h2f_axi_master_arid
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                 // hps_0:h2f_ARLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_arlock
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                 // hps_0:h2f_AWLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_awlock
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                 // hps_0:h2f_AWADDR -> mm_interconnect_1:hps_0_h2f_axi_master_awaddr
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                  // mm_interconnect_1:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire          hps_0_h2f_axi_master_arready;                                // mm_interconnect_1:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire   [63:0] hps_0_h2f_axi_master_rdata;                                  // mm_interconnect_1:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire          hps_0_h2f_axi_master_awready;                                // mm_interconnect_1:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                // hps_0:h2f_ARBURST -> mm_interconnect_1:hps_0_h2f_axi_master_arburst
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                 // hps_0:h2f_ARSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_arsize
	wire          hps_0_h2f_axi_master_bready;                                 // hps_0:h2f_BREADY -> mm_interconnect_1:hps_0_h2f_axi_master_bready
	wire          hps_0_h2f_axi_master_rlast;                                  // mm_interconnect_1:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire          hps_0_h2f_axi_master_wlast;                                  // hps_0:h2f_WLAST -> mm_interconnect_1:hps_0_h2f_axi_master_wlast
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                  // mm_interconnect_1:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire   [11:0] hps_0_h2f_axi_master_awid;                                   // hps_0:h2f_AWID -> mm_interconnect_1:hps_0_h2f_axi_master_awid
	wire   [11:0] hps_0_h2f_axi_master_bid;                                    // mm_interconnect_1:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire          hps_0_h2f_axi_master_bvalid;                                 // mm_interconnect_1:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                 // hps_0:h2f_AWSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_awsize
	wire          hps_0_h2f_axi_master_awvalid;                                // hps_0:h2f_AWVALID -> mm_interconnect_1:hps_0_h2f_axi_master_awvalid
	wire          hps_0_h2f_axi_master_rvalid;                                 // mm_interconnect_1:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire          mm_interconnect_1_sdram_controller_s1_chipselect;            // mm_interconnect_1:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire   [15:0] mm_interconnect_1_sdram_controller_s1_readdata;              // sdram_controller:za_data -> mm_interconnect_1:sdram_controller_s1_readdata
	wire          mm_interconnect_1_sdram_controller_s1_waitrequest;           // sdram_controller:za_waitrequest -> mm_interconnect_1:sdram_controller_s1_waitrequest
	wire   [24:0] mm_interconnect_1_sdram_controller_s1_address;               // mm_interconnect_1:sdram_controller_s1_address -> sdram_controller:az_addr
	wire          mm_interconnect_1_sdram_controller_s1_read;                  // mm_interconnect_1:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire    [1:0] mm_interconnect_1_sdram_controller_s1_byteenable;            // mm_interconnect_1:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire          mm_interconnect_1_sdram_controller_s1_readdatavalid;         // sdram_controller:za_valid -> mm_interconnect_1:sdram_controller_s1_readdatavalid
	wire          mm_interconnect_1_sdram_controller_s1_write;                 // mm_interconnect_1:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire   [15:0] mm_interconnect_1_sdram_controller_s1_writedata;             // mm_interconnect_1:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                             // hps_0:h2f_lw_AWBURST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awburst
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                               // hps_0:h2f_lw_ARLEN -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arlen
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                               // hps_0:h2f_lw_WSTRB -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_wready;                              // mm_interconnect_2:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                                 // mm_interconnect_2:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_rready;                              // hps_0:h2f_lw_RREADY -> mm_interconnect_2:hps_0_h2f_lw_axi_master_rready
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                               // hps_0:h2f_lw_AWLEN -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awlen
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                                 // hps_0:h2f_lw_WID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wid
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                             // hps_0:h2f_lw_ARCACHE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arcache
	wire          hps_0_h2f_lw_axi_master_wvalid;                              // hps_0:h2f_lw_WVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                              // hps_0:h2f_lw_ARADDR -> mm_interconnect_2:hps_0_h2f_lw_axi_master_araddr
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                              // hps_0:h2f_lw_ARPROT -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arprot
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                              // hps_0:h2f_lw_AWPROT -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awprot
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                               // hps_0:h2f_lw_WDATA -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_arvalid;                             // hps_0:h2f_lw_ARVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                             // hps_0:h2f_lw_AWCACHE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awcache
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                                // hps_0:h2f_lw_ARID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arid
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                              // hps_0:h2f_lw_ARLOCK -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                              // hps_0:h2f_lw_AWLOCK -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awlock
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                              // hps_0:h2f_lw_AWADDR -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                               // mm_interconnect_2:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire          hps_0_h2f_lw_axi_master_arready;                             // mm_interconnect_2:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                               // mm_interconnect_2:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire          hps_0_h2f_lw_axi_master_awready;                             // mm_interconnect_2:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                             // hps_0:h2f_lw_ARBURST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arburst
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                              // hps_0:h2f_lw_ARSIZE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arsize
	wire          hps_0_h2f_lw_axi_master_bready;                              // hps_0:h2f_lw_BREADY -> mm_interconnect_2:hps_0_h2f_lw_axi_master_bready
	wire          hps_0_h2f_lw_axi_master_rlast;                               // mm_interconnect_2:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire          hps_0_h2f_lw_axi_master_wlast;                               // hps_0:h2f_lw_WLAST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wlast
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                               // mm_interconnect_2:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                                // hps_0:h2f_lw_AWID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awid
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                                 // mm_interconnect_2:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire          hps_0_h2f_lw_axi_master_bvalid;                              // mm_interconnect_2:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                              // hps_0:h2f_lw_AWSIZE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awsize
	wire          hps_0_h2f_lw_axi_master_awvalid;                             // hps_0:h2f_lw_AWVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awvalid
	wire          hps_0_h2f_lw_axi_master_rvalid;                              // mm_interconnect_2:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire          mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire   [31:0] mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_readdata
	wire          mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire          mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire          mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire   [31:0] mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [31:0] mm_interconnect_2_alt_vip_vfr_0_avalon_slave_readdata;       // alt_vip_vfr_0:slave_readdata -> mm_interconnect_2:alt_vip_vfr_0_avalon_slave_readdata
	wire    [4:0] mm_interconnect_2_alt_vip_vfr_0_avalon_slave_address;        // mm_interconnect_2:alt_vip_vfr_0_avalon_slave_address -> alt_vip_vfr_0:slave_address
	wire          mm_interconnect_2_alt_vip_vfr_0_avalon_slave_read;           // mm_interconnect_2:alt_vip_vfr_0_avalon_slave_read -> alt_vip_vfr_0:slave_read
	wire          mm_interconnect_2_alt_vip_vfr_0_avalon_slave_write;          // mm_interconnect_2:alt_vip_vfr_0_avalon_slave_write -> alt_vip_vfr_0:slave_write
	wire   [31:0] mm_interconnect_2_alt_vip_vfr_0_avalon_slave_writedata;      // mm_interconnect_2:alt_vip_vfr_0_avalon_slave_writedata -> alt_vip_vfr_0:slave_writedata
	wire   [31:0] mm_interconnect_2_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_2:sysid_qsys_0_control_slave_readdata
	wire    [0:0] mm_interconnect_2_sysid_qsys_0_control_slave_address;        // mm_interconnect_2:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire   [31:0] mm_interconnect_2_switches_s1_readdata;                      // switches:readdata -> mm_interconnect_2:switches_s1_readdata
	wire    [1:0] mm_interconnect_2_switches_s1_address;                       // mm_interconnect_2:switches_s1_address -> switches:address
	wire          mm_interconnect_2_led_s1_chipselect;                         // mm_interconnect_2:led_s1_chipselect -> led:chipselect
	wire   [31:0] mm_interconnect_2_led_s1_readdata;                           // led:readdata -> mm_interconnect_2:led_s1_readdata
	wire    [1:0] mm_interconnect_2_led_s1_address;                            // mm_interconnect_2:led_s1_address -> led:address
	wire          mm_interconnect_2_led_s1_write;                              // mm_interconnect_2:led_s1_write -> led:write_n
	wire   [31:0] mm_interconnect_2_led_s1_writedata;                          // mm_interconnect_2:led_s1_writedata -> led:writedata
	wire          mm_interconnect_2_donesignal_s1_chipselect;                  // mm_interconnect_2:doneSignal_s1_chipselect -> doneSignal:chipselect
	wire   [31:0] mm_interconnect_2_donesignal_s1_readdata;                    // doneSignal:readdata -> mm_interconnect_2:doneSignal_s1_readdata
	wire    [1:0] mm_interconnect_2_donesignal_s1_address;                     // mm_interconnect_2:doneSignal_s1_address -> doneSignal:address
	wire          mm_interconnect_2_donesignal_s1_write;                       // mm_interconnect_2:doneSignal_s1_write -> doneSignal:write_n
	wire   [31:0] mm_interconnect_2_donesignal_s1_writedata;                   // mm_interconnect_2:doneSignal_s1_writedata -> doneSignal:writedata
	wire          mm_interconnect_2_startsignal_s1_chipselect;                 // mm_interconnect_2:startSignal_s1_chipselect -> startSignal:chipselect
	wire   [31:0] mm_interconnect_2_startsignal_s1_readdata;                   // startSignal:readdata -> mm_interconnect_2:startSignal_s1_readdata
	wire    [1:0] mm_interconnect_2_startsignal_s1_address;                    // mm_interconnect_2:startSignal_s1_address -> startSignal:address
	wire          mm_interconnect_2_startsignal_s1_write;                      // mm_interconnect_2:startSignal_s1_write -> startSignal:write_n
	wire   [31:0] mm_interconnect_2_startsignal_s1_writedata;                  // mm_interconnect_2:startSignal_s1_writedata -> startSignal:writedata
	wire          irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire   [31:0] hps_0_f2h_irq0_irq;                                          // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                          // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [alt_vip_itc_0:rst, alt_vip_vfr_0:reset, mm_interconnect_2:alt_vip_vfr_0_clock_reset_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [alt_vip_vfr_0:master_reset, doneSignal:reset_n, jtag_uart_0:rst_n, led:reset_n, mm_interconnect_0:alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset_reset, mm_interconnect_1:sdram_master_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:jtag_uart_0_reset_reset_bridge_in_reset_reset, sdram_controller:reset_n, sdram_master_0:reset_n, startSignal:reset_n, switches:reset_n, sysid_qsys_0:reset_n]
	wire          rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [mm_interconnect_0:hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]

	alt_vipitc131_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (4),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (1024),
		.V_ACTIVE_LINES                (768),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (1920),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (1919),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (136),
		.H_FRONT_PORCH                 (24),
		.H_BACK_PORCH                  (160),
		.V_SYNC_LENGTH                 (6),
		.V_FRONT_PORCH                 (3),
		.V_BACK_PORCH                  (29),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_0 (
		.is_clk        (pll_0_outclk0_clk),                                   //       is_clk_rst.clk
		.rst           (rst_controller_reset_out_reset),                      // is_clk_rst_reset.reset
		.is_data       (alt_vip_vfr_0_avalon_streaming_source_data),          //              din.data
		.is_valid      (alt_vip_vfr_0_avalon_streaming_source_valid),         //                 .valid
		.is_ready      (alt_vip_vfr_0_avalon_streaming_source_ready),         //                 .ready
		.is_sop        (alt_vip_vfr_0_avalon_streaming_source_startofpacket), //                 .startofpacket
		.is_eop        (alt_vip_vfr_0_avalon_streaming_source_endofpacket),   //                 .endofpacket
		.vid_clk       (alt_vip_itc_0_clocked_video_vid_clk),                 //    clocked_video.export
		.vid_data      (alt_vip_itc_0_clocked_video_vid_data),                //                 .export
		.underflow     (alt_vip_itc_0_clocked_video_underflow),               //                 .export
		.vid_datavalid (alt_vip_itc_0_clocked_video_vid_datavalid),           //                 .export
		.vid_v_sync    (alt_vip_itc_0_clocked_video_vid_v_sync),              //                 .export
		.vid_h_sync    (alt_vip_itc_0_clocked_video_vid_h_sync),              //                 .export
		.vid_f         (alt_vip_itc_0_clocked_video_vid_f),                   //                 .export
		.vid_h         (alt_vip_itc_0_clocked_video_vid_h),                   //                 .export
		.vid_v         (alt_vip_itc_0_clocked_video_vid_v)                    //                 .export
	);

	alt_vipvfr131_vfr #(
		.BITS_PER_PIXEL_PER_COLOR_PLANE (8),
		.NUMBER_OF_CHANNELS_IN_PARALLEL (4),
		.NUMBER_OF_CHANNELS_IN_SEQUENCE (1),
		.MAX_IMAGE_WIDTH                (1024),
		.MAX_IMAGE_HEIGHT               (768),
		.MEM_PORT_WIDTH                 (128),
		.RMASTER_FIFO_DEPTH             (64),
		.RMASTER_BURST_TARGET           (32),
		.CLOCKS_ARE_SEPARATE            (1)
	) alt_vip_vfr_0 (
		.clock                (pll_0_outclk0_clk),                                      //             clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                         //       clock_reset_reset.reset
		.master_clock         (sys_clk_sys_clk_clk),                                    //            clock_master.clk
		.master_reset         (rst_controller_001_reset_out_reset),                     //      clock_master_reset.reset
		.slave_address        (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_address),   //            avalon_slave.address
		.slave_write          (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_write),     //                        .write
		.slave_writedata      (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_writedata), //                        .writedata
		.slave_read           (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_read),      //                        .read
		.slave_readdata       (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_readdata),  //                        .readdata
		.slave_irq            (),                                                       //        interrupt_sender.irq
		.dout_data            (alt_vip_vfr_0_avalon_streaming_source_data),             // avalon_streaming_source.data
		.dout_valid           (alt_vip_vfr_0_avalon_streaming_source_valid),            //                        .valid
		.dout_ready           (alt_vip_vfr_0_avalon_streaming_source_ready),            //                        .ready
		.dout_startofpacket   (alt_vip_vfr_0_avalon_streaming_source_startofpacket),    //                        .startofpacket
		.dout_endofpacket     (alt_vip_vfr_0_avalon_streaming_source_endofpacket),      //                        .endofpacket
		.master_address       (alt_vip_vfr_0_avalon_master_address),                    //           avalon_master.address
		.master_burstcount    (alt_vip_vfr_0_avalon_master_burstcount),                 //                        .burstcount
		.master_readdata      (alt_vip_vfr_0_avalon_master_readdata),                   //                        .readdata
		.master_read          (alt_vip_vfr_0_avalon_master_read),                       //                        .read
		.master_readdatavalid (alt_vip_vfr_0_avalon_master_readdatavalid),              //                        .readdatavalid
		.master_waitrequest   (alt_vip_vfr_0_avalon_master_waitrequest)                 //                        .waitrequest
	);

	mysystem_doneSignal donesignal (
		.clk        (sys_clk_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_2_donesignal_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_donesignal_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_donesignal_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_donesignal_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_donesignal_s1_readdata),   //                    .readdata
		.in_port    (donesig_export)                              // external_connection.export
	);

	mysystem_hps_0 #(
		.F2S_Width (3),
		.S2F_Width (2)
	) hps_0 (
		.f2h_boot_from_fpga_ready      (),                                              // f2h_boot_from_fpga.boot_from_fpga_ready
		.f2h_boot_from_fpga_on_failure (),                                              //                   .boot_from_fpga_on_failure
		.mem_a                         (memory_mem_a),                                  //             memory.mem_a
		.mem_ba                        (memory_mem_ba),                                 //                   .mem_ba
		.mem_ck                        (memory_mem_ck),                                 //                   .mem_ck
		.mem_ck_n                      (memory_mem_ck_n),                               //                   .mem_ck_n
		.mem_cke                       (memory_mem_cke),                                //                   .mem_cke
		.mem_cs_n                      (memory_mem_cs_n),                               //                   .mem_cs_n
		.mem_ras_n                     (memory_mem_ras_n),                              //                   .mem_ras_n
		.mem_cas_n                     (memory_mem_cas_n),                              //                   .mem_cas_n
		.mem_we_n                      (memory_mem_we_n),                               //                   .mem_we_n
		.mem_reset_n                   (memory_mem_reset_n),                            //                   .mem_reset_n
		.mem_dq                        (memory_mem_dq),                                 //                   .mem_dq
		.mem_dqs                       (memory_mem_dqs),                                //                   .mem_dqs
		.mem_dqs_n                     (memory_mem_dqs_n),                              //                   .mem_dqs_n
		.mem_odt                       (memory_mem_odt),                                //                   .mem_odt
		.mem_dm                        (memory_mem_dm),                                 //                   .mem_dm
		.oct_rzqin                     (memory_oct_rzqin),                              //                   .oct_rzqin
		.hps_io_sdio_inst_CMD          (hps_io_hps_io_sdio_inst_CMD),                   //             hps_io.hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0           (hps_io_hps_io_sdio_inst_D0),                    //                   .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1           (hps_io_hps_io_sdio_inst_D1),                    //                   .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK          (hps_io_hps_io_sdio_inst_CLK),                   //                   .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2           (hps_io_hps_io_sdio_inst_D2),                    //                   .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3           (hps_io_hps_io_sdio_inst_D3),                    //                   .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0           (hps_io_hps_io_usb1_inst_D0),                    //                   .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1           (hps_io_hps_io_usb1_inst_D1),                    //                   .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2           (hps_io_hps_io_usb1_inst_D2),                    //                   .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3           (hps_io_hps_io_usb1_inst_D3),                    //                   .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4           (hps_io_hps_io_usb1_inst_D4),                    //                   .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5           (hps_io_hps_io_usb1_inst_D5),                    //                   .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6           (hps_io_hps_io_usb1_inst_D6),                    //                   .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7           (hps_io_hps_io_usb1_inst_D7),                    //                   .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK          (hps_io_hps_io_usb1_inst_CLK),                   //                   .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP          (hps_io_hps_io_usb1_inst_STP),                   //                   .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR          (hps_io_hps_io_usb1_inst_DIR),                   //                   .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT          (hps_io_hps_io_usb1_inst_NXT),                   //                   .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX          (hps_io_hps_io_uart0_inst_RX),                   //                   .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX          (hps_io_hps_io_uart0_inst_TX),                   //                   .hps_io_uart0_inst_TX
		.h2f_rst_n                     (hps_0_h2f_reset_reset_n),                       //          h2f_reset.reset_n
		.h2f_axi_clk                   (sys_clk_sys_clk_clk),                           //      h2f_axi_clock.clk
		.h2f_AWID                      (hps_0_h2f_axi_master_awid),                     //     h2f_axi_master.awid
		.h2f_AWADDR                    (hps_0_h2f_axi_master_awaddr),                   //                   .awaddr
		.h2f_AWLEN                     (hps_0_h2f_axi_master_awlen),                    //                   .awlen
		.h2f_AWSIZE                    (hps_0_h2f_axi_master_awsize),                   //                   .awsize
		.h2f_AWBURST                   (hps_0_h2f_axi_master_awburst),                  //                   .awburst
		.h2f_AWLOCK                    (hps_0_h2f_axi_master_awlock),                   //                   .awlock
		.h2f_AWCACHE                   (hps_0_h2f_axi_master_awcache),                  //                   .awcache
		.h2f_AWPROT                    (hps_0_h2f_axi_master_awprot),                   //                   .awprot
		.h2f_AWVALID                   (hps_0_h2f_axi_master_awvalid),                  //                   .awvalid
		.h2f_AWREADY                   (hps_0_h2f_axi_master_awready),                  //                   .awready
		.h2f_WID                       (hps_0_h2f_axi_master_wid),                      //                   .wid
		.h2f_WDATA                     (hps_0_h2f_axi_master_wdata),                    //                   .wdata
		.h2f_WSTRB                     (hps_0_h2f_axi_master_wstrb),                    //                   .wstrb
		.h2f_WLAST                     (hps_0_h2f_axi_master_wlast),                    //                   .wlast
		.h2f_WVALID                    (hps_0_h2f_axi_master_wvalid),                   //                   .wvalid
		.h2f_WREADY                    (hps_0_h2f_axi_master_wready),                   //                   .wready
		.h2f_BID                       (hps_0_h2f_axi_master_bid),                      //                   .bid
		.h2f_BRESP                     (hps_0_h2f_axi_master_bresp),                    //                   .bresp
		.h2f_BVALID                    (hps_0_h2f_axi_master_bvalid),                   //                   .bvalid
		.h2f_BREADY                    (hps_0_h2f_axi_master_bready),                   //                   .bready
		.h2f_ARID                      (hps_0_h2f_axi_master_arid),                     //                   .arid
		.h2f_ARADDR                    (hps_0_h2f_axi_master_araddr),                   //                   .araddr
		.h2f_ARLEN                     (hps_0_h2f_axi_master_arlen),                    //                   .arlen
		.h2f_ARSIZE                    (hps_0_h2f_axi_master_arsize),                   //                   .arsize
		.h2f_ARBURST                   (hps_0_h2f_axi_master_arburst),                  //                   .arburst
		.h2f_ARLOCK                    (hps_0_h2f_axi_master_arlock),                   //                   .arlock
		.h2f_ARCACHE                   (hps_0_h2f_axi_master_arcache),                  //                   .arcache
		.h2f_ARPROT                    (hps_0_h2f_axi_master_arprot),                   //                   .arprot
		.h2f_ARVALID                   (hps_0_h2f_axi_master_arvalid),                  //                   .arvalid
		.h2f_ARREADY                   (hps_0_h2f_axi_master_arready),                  //                   .arready
		.h2f_RID                       (hps_0_h2f_axi_master_rid),                      //                   .rid
		.h2f_RDATA                     (hps_0_h2f_axi_master_rdata),                    //                   .rdata
		.h2f_RRESP                     (hps_0_h2f_axi_master_rresp),                    //                   .rresp
		.h2f_RLAST                     (hps_0_h2f_axi_master_rlast),                    //                   .rlast
		.h2f_RVALID                    (hps_0_h2f_axi_master_rvalid),                   //                   .rvalid
		.h2f_RREADY                    (hps_0_h2f_axi_master_rready),                   //                   .rready
		.f2h_axi_clk                   (sys_clk_sys_clk_clk),                           //      f2h_axi_clock.clk
		.f2h_AWID                      (mm_interconnect_0_hps_0_f2h_axi_slave_awid),    //      f2h_axi_slave.awid
		.f2h_AWADDR                    (mm_interconnect_0_hps_0_f2h_axi_slave_awaddr),  //                   .awaddr
		.f2h_AWLEN                     (mm_interconnect_0_hps_0_f2h_axi_slave_awlen),   //                   .awlen
		.f2h_AWSIZE                    (mm_interconnect_0_hps_0_f2h_axi_slave_awsize),  //                   .awsize
		.f2h_AWBURST                   (mm_interconnect_0_hps_0_f2h_axi_slave_awburst), //                   .awburst
		.f2h_AWLOCK                    (mm_interconnect_0_hps_0_f2h_axi_slave_awlock),  //                   .awlock
		.f2h_AWCACHE                   (mm_interconnect_0_hps_0_f2h_axi_slave_awcache), //                   .awcache
		.f2h_AWPROT                    (mm_interconnect_0_hps_0_f2h_axi_slave_awprot),  //                   .awprot
		.f2h_AWVALID                   (mm_interconnect_0_hps_0_f2h_axi_slave_awvalid), //                   .awvalid
		.f2h_AWREADY                   (mm_interconnect_0_hps_0_f2h_axi_slave_awready), //                   .awready
		.f2h_AWUSER                    (mm_interconnect_0_hps_0_f2h_axi_slave_awuser),  //                   .awuser
		.f2h_WID                       (mm_interconnect_0_hps_0_f2h_axi_slave_wid),     //                   .wid
		.f2h_WDATA                     (mm_interconnect_0_hps_0_f2h_axi_slave_wdata),   //                   .wdata
		.f2h_WSTRB                     (mm_interconnect_0_hps_0_f2h_axi_slave_wstrb),   //                   .wstrb
		.f2h_WLAST                     (mm_interconnect_0_hps_0_f2h_axi_slave_wlast),   //                   .wlast
		.f2h_WVALID                    (mm_interconnect_0_hps_0_f2h_axi_slave_wvalid),  //                   .wvalid
		.f2h_WREADY                    (mm_interconnect_0_hps_0_f2h_axi_slave_wready),  //                   .wready
		.f2h_BID                       (mm_interconnect_0_hps_0_f2h_axi_slave_bid),     //                   .bid
		.f2h_BRESP                     (mm_interconnect_0_hps_0_f2h_axi_slave_bresp),   //                   .bresp
		.f2h_BVALID                    (mm_interconnect_0_hps_0_f2h_axi_slave_bvalid),  //                   .bvalid
		.f2h_BREADY                    (mm_interconnect_0_hps_0_f2h_axi_slave_bready),  //                   .bready
		.f2h_ARID                      (mm_interconnect_0_hps_0_f2h_axi_slave_arid),    //                   .arid
		.f2h_ARADDR                    (mm_interconnect_0_hps_0_f2h_axi_slave_araddr),  //                   .araddr
		.f2h_ARLEN                     (mm_interconnect_0_hps_0_f2h_axi_slave_arlen),   //                   .arlen
		.f2h_ARSIZE                    (mm_interconnect_0_hps_0_f2h_axi_slave_arsize),  //                   .arsize
		.f2h_ARBURST                   (mm_interconnect_0_hps_0_f2h_axi_slave_arburst), //                   .arburst
		.f2h_ARLOCK                    (mm_interconnect_0_hps_0_f2h_axi_slave_arlock),  //                   .arlock
		.f2h_ARCACHE                   (mm_interconnect_0_hps_0_f2h_axi_slave_arcache), //                   .arcache
		.f2h_ARPROT                    (mm_interconnect_0_hps_0_f2h_axi_slave_arprot),  //                   .arprot
		.f2h_ARVALID                   (mm_interconnect_0_hps_0_f2h_axi_slave_arvalid), //                   .arvalid
		.f2h_ARREADY                   (mm_interconnect_0_hps_0_f2h_axi_slave_arready), //                   .arready
		.f2h_ARUSER                    (mm_interconnect_0_hps_0_f2h_axi_slave_aruser),  //                   .aruser
		.f2h_RID                       (mm_interconnect_0_hps_0_f2h_axi_slave_rid),     //                   .rid
		.f2h_RDATA                     (mm_interconnect_0_hps_0_f2h_axi_slave_rdata),   //                   .rdata
		.f2h_RRESP                     (mm_interconnect_0_hps_0_f2h_axi_slave_rresp),   //                   .rresp
		.f2h_RLAST                     (mm_interconnect_0_hps_0_f2h_axi_slave_rlast),   //                   .rlast
		.f2h_RVALID                    (mm_interconnect_0_hps_0_f2h_axi_slave_rvalid),  //                   .rvalid
		.f2h_RREADY                    (mm_interconnect_0_hps_0_f2h_axi_slave_rready),  //                   .rready
		.h2f_lw_axi_clk                (sys_clk_sys_clk_clk),                           //   h2f_lw_axi_clock.clk
		.h2f_lw_AWID                   (hps_0_h2f_lw_axi_master_awid),                  //  h2f_lw_axi_master.awid
		.h2f_lw_AWADDR                 (hps_0_h2f_lw_axi_master_awaddr),                //                   .awaddr
		.h2f_lw_AWLEN                  (hps_0_h2f_lw_axi_master_awlen),                 //                   .awlen
		.h2f_lw_AWSIZE                 (hps_0_h2f_lw_axi_master_awsize),                //                   .awsize
		.h2f_lw_AWBURST                (hps_0_h2f_lw_axi_master_awburst),               //                   .awburst
		.h2f_lw_AWLOCK                 (hps_0_h2f_lw_axi_master_awlock),                //                   .awlock
		.h2f_lw_AWCACHE                (hps_0_h2f_lw_axi_master_awcache),               //                   .awcache
		.h2f_lw_AWPROT                 (hps_0_h2f_lw_axi_master_awprot),                //                   .awprot
		.h2f_lw_AWVALID                (hps_0_h2f_lw_axi_master_awvalid),               //                   .awvalid
		.h2f_lw_AWREADY                (hps_0_h2f_lw_axi_master_awready),               //                   .awready
		.h2f_lw_WID                    (hps_0_h2f_lw_axi_master_wid),                   //                   .wid
		.h2f_lw_WDATA                  (hps_0_h2f_lw_axi_master_wdata),                 //                   .wdata
		.h2f_lw_WSTRB                  (hps_0_h2f_lw_axi_master_wstrb),                 //                   .wstrb
		.h2f_lw_WLAST                  (hps_0_h2f_lw_axi_master_wlast),                 //                   .wlast
		.h2f_lw_WVALID                 (hps_0_h2f_lw_axi_master_wvalid),                //                   .wvalid
		.h2f_lw_WREADY                 (hps_0_h2f_lw_axi_master_wready),                //                   .wready
		.h2f_lw_BID                    (hps_0_h2f_lw_axi_master_bid),                   //                   .bid
		.h2f_lw_BRESP                  (hps_0_h2f_lw_axi_master_bresp),                 //                   .bresp
		.h2f_lw_BVALID                 (hps_0_h2f_lw_axi_master_bvalid),                //                   .bvalid
		.h2f_lw_BREADY                 (hps_0_h2f_lw_axi_master_bready),                //                   .bready
		.h2f_lw_ARID                   (hps_0_h2f_lw_axi_master_arid),                  //                   .arid
		.h2f_lw_ARADDR                 (hps_0_h2f_lw_axi_master_araddr),                //                   .araddr
		.h2f_lw_ARLEN                  (hps_0_h2f_lw_axi_master_arlen),                 //                   .arlen
		.h2f_lw_ARSIZE                 (hps_0_h2f_lw_axi_master_arsize),                //                   .arsize
		.h2f_lw_ARBURST                (hps_0_h2f_lw_axi_master_arburst),               //                   .arburst
		.h2f_lw_ARLOCK                 (hps_0_h2f_lw_axi_master_arlock),                //                   .arlock
		.h2f_lw_ARCACHE                (hps_0_h2f_lw_axi_master_arcache),               //                   .arcache
		.h2f_lw_ARPROT                 (hps_0_h2f_lw_axi_master_arprot),                //                   .arprot
		.h2f_lw_ARVALID                (hps_0_h2f_lw_axi_master_arvalid),               //                   .arvalid
		.h2f_lw_ARREADY                (hps_0_h2f_lw_axi_master_arready),               //                   .arready
		.h2f_lw_RID                    (hps_0_h2f_lw_axi_master_rid),                   //                   .rid
		.h2f_lw_RDATA                  (hps_0_h2f_lw_axi_master_rdata),                 //                   .rdata
		.h2f_lw_RRESP                  (hps_0_h2f_lw_axi_master_rresp),                 //                   .rresp
		.h2f_lw_RLAST                  (hps_0_h2f_lw_axi_master_rlast),                 //                   .rlast
		.h2f_lw_RVALID                 (hps_0_h2f_lw_axi_master_rvalid),                //                   .rvalid
		.h2f_lw_RREADY                 (hps_0_h2f_lw_axi_master_rready),                //                   .rready
		.f2h_irq_p0                    (hps_0_f2h_irq0_irq),                            //           f2h_irq0.irq
		.f2h_irq_p1                    (hps_0_f2h_irq1_irq)                             //           f2h_irq1.irq
	);

	mysystem_jtag_uart_0 jtag_uart_0 (
		.clk            (sys_clk_sys_clk_clk),                                         //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	mysystem_led led (
		.clk        (sys_clk_sys_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_2_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	mysystem_pll_0 pll_0 (
		.refclk   (sys_clk_sys_clk_clk),        //  refclk.clk
		.rst      (sys_clk_reset_source_reset), //   reset.reset
		.outclk_0 (pll_0_outclk0_clk),          // outclk0.clk
		.locked   ()                            //  locked.export
	);

	mysystem_pll_1 pll_1 (
		.refclk   (sys_clk_sys_clk_clk),        //  refclk.clk
		.rst      (sys_clk_reset_source_reset), //   reset.reset
		.outclk_0 (clk_65_clk),                 // outclk0.clk
		.locked   ()                            //  locked.export
	);

	mysystem_sdram_controller sdram_controller (
		.clk            (sys_clk_sys_clk_clk),                                 //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                 // reset.reset_n
		.az_addr        (mm_interconnect_1_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_1_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_1_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_1_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_1_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_1_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_1_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_1_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_1_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                     //  wire.export
		.zs_ba          (sdram_wire_ba),                                       //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                    //      .export
		.zs_cke         (sdram_wire_cke),                                      //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                     //      .export
		.zs_dq          (sdram_wire_dq),                                       //      .export
		.zs_dqm         (sdram_wire_dqm),                                      //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                    //      .export
		.zs_we_n        (sdram_wire_we_n)                                      //      .export
	);

	sdram_master sdram_master_0 (
		.clk           (sys_clk_sys_clk_clk),                        //         clock.clk
		.reset_n       (~rst_controller_001_reset_out_reset),        //         reset.reset_n
		.read_n        (sdram_master_0_avalon_master_read),          // avalon_master.read_n
		.write_n       (sdram_master_0_avalon_master_write),         //              .write_n
		.chipselect    (sdram_master_0_avalon_master_chipselect),    //              .chipselect
		.waitrequest   (sdram_master_0_avalon_master_waitrequest),   //              .waitrequest
		.address       (sdram_master_0_avalon_master_address),       //              .address
		.byteenable    (sdram_master_0_avalon_master_byteenable),    //              .byteenable
		.readdatavalid (sdram_master_0_avalon_master_readdatavalid), //              .readdatavalid
		.readdata      (sdram_master_0_avalon_master_readdata),      //              .readdata
		.writedata     (sdram_master_0_avalon_master_writedata),     //              .writedata
		.s             (sdramstartstop_readdata),                    //   conduit_end.readdata
		.startSig      (sdramstartstop_beginbursttransfer),          //              .beginbursttransfer
		.doneSig       (sdramstartstop_writeresponsevalid_n)         //              .writeresponsevalid_n
	);

	mysystem_startSignal startsignal (
		.clk        (sys_clk_sys_clk_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_2_startsignal_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_startsignal_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_startsignal_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_startsignal_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_startsignal_s1_readdata),   //                    .readdata
		.out_port   (startsig_export)                              // external_connection.export
	);

	mysystem_switches switches (
		.clk      (sys_clk_sys_clk_clk),                    //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_2_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_switches_s1_readdata), //                    .readdata
		.in_port  (switches_external_connection_export)     // external_connection.export
	);

	mysystem_sys_clk sys_clk (
		.ref_clk_clk        (system_ref_clk_clk),         //      ref_clk.clk
		.ref_reset_reset    (system_ref_reset_reset),     //    ref_reset.reset
		.sys_clk_clk        (sys_clk_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),              //    sdram_clk.clk
		.reset_source_reset (sys_clk_reset_source_reset)  // reset_source.reset
	);

	mysystem_sysid_qsys_0 sysid_qsys_0 (
		.clock    (sys_clk_sys_clk_clk),                                   //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_2_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_2_sysid_qsys_0_control_slave_address)   //              .address
	);

	mysystem_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_f2h_axi_slave_awid                                         (mm_interconnect_0_hps_0_f2h_axi_slave_awid),    //                                        hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awaddr),  //                                                           .awaddr
		.hps_0_f2h_axi_slave_awlen                                        (mm_interconnect_0_hps_0_f2h_axi_slave_awlen),   //                                                           .awlen
		.hps_0_f2h_axi_slave_awsize                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awsize),  //                                                           .awsize
		.hps_0_f2h_axi_slave_awburst                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awburst), //                                                           .awburst
		.hps_0_f2h_axi_slave_awlock                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awlock),  //                                                           .awlock
		.hps_0_f2h_axi_slave_awcache                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awcache), //                                                           .awcache
		.hps_0_f2h_axi_slave_awprot                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awprot),  //                                                           .awprot
		.hps_0_f2h_axi_slave_awuser                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awuser),  //                                                           .awuser
		.hps_0_f2h_axi_slave_awvalid                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awvalid), //                                                           .awvalid
		.hps_0_f2h_axi_slave_awready                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awready), //                                                           .awready
		.hps_0_f2h_axi_slave_wid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_wid),     //                                                           .wid
		.hps_0_f2h_axi_slave_wdata                                        (mm_interconnect_0_hps_0_f2h_axi_slave_wdata),   //                                                           .wdata
		.hps_0_f2h_axi_slave_wstrb                                        (mm_interconnect_0_hps_0_f2h_axi_slave_wstrb),   //                                                           .wstrb
		.hps_0_f2h_axi_slave_wlast                                        (mm_interconnect_0_hps_0_f2h_axi_slave_wlast),   //                                                           .wlast
		.hps_0_f2h_axi_slave_wvalid                                       (mm_interconnect_0_hps_0_f2h_axi_slave_wvalid),  //                                                           .wvalid
		.hps_0_f2h_axi_slave_wready                                       (mm_interconnect_0_hps_0_f2h_axi_slave_wready),  //                                                           .wready
		.hps_0_f2h_axi_slave_bid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_bid),     //                                                           .bid
		.hps_0_f2h_axi_slave_bresp                                        (mm_interconnect_0_hps_0_f2h_axi_slave_bresp),   //                                                           .bresp
		.hps_0_f2h_axi_slave_bvalid                                       (mm_interconnect_0_hps_0_f2h_axi_slave_bvalid),  //                                                           .bvalid
		.hps_0_f2h_axi_slave_bready                                       (mm_interconnect_0_hps_0_f2h_axi_slave_bready),  //                                                           .bready
		.hps_0_f2h_axi_slave_arid                                         (mm_interconnect_0_hps_0_f2h_axi_slave_arid),    //                                                           .arid
		.hps_0_f2h_axi_slave_araddr                                       (mm_interconnect_0_hps_0_f2h_axi_slave_araddr),  //                                                           .araddr
		.hps_0_f2h_axi_slave_arlen                                        (mm_interconnect_0_hps_0_f2h_axi_slave_arlen),   //                                                           .arlen
		.hps_0_f2h_axi_slave_arsize                                       (mm_interconnect_0_hps_0_f2h_axi_slave_arsize),  //                                                           .arsize
		.hps_0_f2h_axi_slave_arburst                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arburst), //                                                           .arburst
		.hps_0_f2h_axi_slave_arlock                                       (mm_interconnect_0_hps_0_f2h_axi_slave_arlock),  //                                                           .arlock
		.hps_0_f2h_axi_slave_arcache                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arcache), //                                                           .arcache
		.hps_0_f2h_axi_slave_arprot                                       (mm_interconnect_0_hps_0_f2h_axi_slave_arprot),  //                                                           .arprot
		.hps_0_f2h_axi_slave_aruser                                       (mm_interconnect_0_hps_0_f2h_axi_slave_aruser),  //                                                           .aruser
		.hps_0_f2h_axi_slave_arvalid                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arvalid), //                                                           .arvalid
		.hps_0_f2h_axi_slave_arready                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arready), //                                                           .arready
		.hps_0_f2h_axi_slave_rid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_rid),     //                                                           .rid
		.hps_0_f2h_axi_slave_rdata                                        (mm_interconnect_0_hps_0_f2h_axi_slave_rdata),   //                                                           .rdata
		.hps_0_f2h_axi_slave_rresp                                        (mm_interconnect_0_hps_0_f2h_axi_slave_rresp),   //                                                           .rresp
		.hps_0_f2h_axi_slave_rlast                                        (mm_interconnect_0_hps_0_f2h_axi_slave_rlast),   //                                                           .rlast
		.hps_0_f2h_axi_slave_rvalid                                       (mm_interconnect_0_hps_0_f2h_axi_slave_rvalid),  //                                                           .rvalid
		.hps_0_f2h_axi_slave_rready                                       (mm_interconnect_0_hps_0_f2h_axi_slave_rready),  //                                                           .rready
		.sys_clk_sys_clk_clk                                              (sys_clk_sys_clk_clk),                           //                                            sys_clk_sys_clk.clk
		.alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),            //     alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset.reset
		.hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),            // hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.alt_vip_vfr_0_avalon_master_address                              (alt_vip_vfr_0_avalon_master_address),           //                                alt_vip_vfr_0_avalon_master.address
		.alt_vip_vfr_0_avalon_master_waitrequest                          (alt_vip_vfr_0_avalon_master_waitrequest),       //                                                           .waitrequest
		.alt_vip_vfr_0_avalon_master_burstcount                           (alt_vip_vfr_0_avalon_master_burstcount),        //                                                           .burstcount
		.alt_vip_vfr_0_avalon_master_read                                 (alt_vip_vfr_0_avalon_master_read),              //                                                           .read
		.alt_vip_vfr_0_avalon_master_readdata                             (alt_vip_vfr_0_avalon_master_readdata),          //                                                           .readdata
		.alt_vip_vfr_0_avalon_master_readdatavalid                        (alt_vip_vfr_0_avalon_master_readdatavalid)      //                                                           .readdatavalid
	);

	mysystem_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                           //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                         //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                          //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                         //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                        //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                         //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                        //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                         //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                        //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                        //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                            //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                          //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                          //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                          //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                         //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                         //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                            //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                          //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                         //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                         //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                           //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                         //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                          //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                         //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                        //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                         //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                        //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                         //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                        //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                        //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                            //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                          //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                          //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                          //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                         //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                         //                                                           .rready
		.sys_clk_sys_clk_clk                                              (sys_clk_sys_clk_clk),                                 //                                            sys_clk_sys_clk.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                  // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.sdram_master_0_reset_reset_bridge_in_reset_reset                 (rst_controller_001_reset_out_reset),                  //                 sdram_master_0_reset_reset_bridge_in_reset.reset
		.sdram_master_0_avalon_master_address                             (sdram_master_0_avalon_master_address),                //                               sdram_master_0_avalon_master.address
		.sdram_master_0_avalon_master_waitrequest                         (sdram_master_0_avalon_master_waitrequest),            //                                                           .waitrequest
		.sdram_master_0_avalon_master_byteenable                          (sdram_master_0_avalon_master_byteenable),             //                                                           .byteenable
		.sdram_master_0_avalon_master_chipselect                          (sdram_master_0_avalon_master_chipselect),             //                                                           .chipselect
		.sdram_master_0_avalon_master_read                                (~sdram_master_0_avalon_master_read),                  //                                                           .read
		.sdram_master_0_avalon_master_readdata                            (sdram_master_0_avalon_master_readdata),               //                                                           .readdata
		.sdram_master_0_avalon_master_readdatavalid                       (sdram_master_0_avalon_master_readdatavalid),          //                                                           .readdatavalid
		.sdram_master_0_avalon_master_write                               (~sdram_master_0_avalon_master_write),                 //                                                           .write
		.sdram_master_0_avalon_master_writedata                           (sdram_master_0_avalon_master_writedata),              //                                                           .writedata
		.sdram_controller_s1_address                                      (mm_interconnect_1_sdram_controller_s1_address),       //                                        sdram_controller_s1.address
		.sdram_controller_s1_write                                        (mm_interconnect_1_sdram_controller_s1_write),         //                                                           .write
		.sdram_controller_s1_read                                         (mm_interconnect_1_sdram_controller_s1_read),          //                                                           .read
		.sdram_controller_s1_readdata                                     (mm_interconnect_1_sdram_controller_s1_readdata),      //                                                           .readdata
		.sdram_controller_s1_writedata                                    (mm_interconnect_1_sdram_controller_s1_writedata),     //                                                           .writedata
		.sdram_controller_s1_byteenable                                   (mm_interconnect_1_sdram_controller_s1_byteenable),    //                                                           .byteenable
		.sdram_controller_s1_readdatavalid                                (mm_interconnect_1_sdram_controller_s1_readdatavalid), //                                                           .readdatavalid
		.sdram_controller_s1_waitrequest                                  (mm_interconnect_1_sdram_controller_s1_waitrequest),   //                                                           .waitrequest
		.sdram_controller_s1_chipselect                                   (mm_interconnect_1_sdram_controller_s1_chipselect)     //                                                           .chipselect
	);

	mysystem_mm_interconnect_2 mm_interconnect_2 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                                //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                              //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                               //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                              //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                             //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                              //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                             //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                              //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                             //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                             //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                                 //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                               //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                               //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                               //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                              //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                              //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                                 //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                               //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                              //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                              //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                                //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                              //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                               //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                              //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                             //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                              //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                             //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                              //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                             //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                             //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                                 //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                               //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                               //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                               //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                              //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                              //                                                              .rready
		.pll_0_outclk0_clk                                                   (pll_0_outclk0_clk),                                           //                                                 pll_0_outclk0.clk
		.sys_clk_sys_clk_clk                                                 (sys_clk_sys_clk_clk),                                         //                                               sys_clk_sys_clk.clk
		.alt_vip_vfr_0_clock_reset_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                              //         alt_vip_vfr_0_clock_reset_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                          // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.jtag_uart_0_reset_reset_bridge_in_reset_reset                       (rst_controller_001_reset_out_reset),                          //                       jtag_uart_0_reset_reset_bridge_in_reset.reset
		.alt_vip_vfr_0_avalon_slave_address                                  (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_address),        //                                    alt_vip_vfr_0_avalon_slave.address
		.alt_vip_vfr_0_avalon_slave_write                                    (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_write),          //                                                              .write
		.alt_vip_vfr_0_avalon_slave_read                                     (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_read),           //                                                              .read
		.alt_vip_vfr_0_avalon_slave_readdata                                 (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_readdata),       //                                                              .readdata
		.alt_vip_vfr_0_avalon_slave_writedata                                (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_writedata),      //                                                              .writedata
		.doneSignal_s1_address                                               (mm_interconnect_2_donesignal_s1_address),                     //                                                 doneSignal_s1.address
		.doneSignal_s1_write                                                 (mm_interconnect_2_donesignal_s1_write),                       //                                                              .write
		.doneSignal_s1_readdata                                              (mm_interconnect_2_donesignal_s1_readdata),                    //                                                              .readdata
		.doneSignal_s1_writedata                                             (mm_interconnect_2_donesignal_s1_writedata),                   //                                                              .writedata
		.doneSignal_s1_chipselect                                            (mm_interconnect_2_donesignal_s1_chipselect),                  //                                                              .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                               (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_address),     //                                 jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                                 (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_write),       //                                                              .write
		.jtag_uart_0_avalon_jtag_slave_read                                  (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_read),        //                                                              .read
		.jtag_uart_0_avalon_jtag_slave_readdata                              (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_readdata),    //                                                              .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                             (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_writedata),   //                                                              .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                           (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                                              .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                            (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                                              .chipselect
		.led_s1_address                                                      (mm_interconnect_2_led_s1_address),                            //                                                        led_s1.address
		.led_s1_write                                                        (mm_interconnect_2_led_s1_write),                              //                                                              .write
		.led_s1_readdata                                                     (mm_interconnect_2_led_s1_readdata),                           //                                                              .readdata
		.led_s1_writedata                                                    (mm_interconnect_2_led_s1_writedata),                          //                                                              .writedata
		.led_s1_chipselect                                                   (mm_interconnect_2_led_s1_chipselect),                         //                                                              .chipselect
		.startSignal_s1_address                                              (mm_interconnect_2_startsignal_s1_address),                    //                                                startSignal_s1.address
		.startSignal_s1_write                                                (mm_interconnect_2_startsignal_s1_write),                      //                                                              .write
		.startSignal_s1_readdata                                             (mm_interconnect_2_startsignal_s1_readdata),                   //                                                              .readdata
		.startSignal_s1_writedata                                            (mm_interconnect_2_startsignal_s1_writedata),                  //                                                              .writedata
		.startSignal_s1_chipselect                                           (mm_interconnect_2_startsignal_s1_chipselect),                 //                                                              .chipselect
		.switches_s1_address                                                 (mm_interconnect_2_switches_s1_address),                       //                                                   switches_s1.address
		.switches_s1_readdata                                                (mm_interconnect_2_switches_s1_readdata),                      //                                                              .readdata
		.sysid_qsys_0_control_slave_address                                  (mm_interconnect_2_sysid_qsys_0_control_slave_address),        //                                    sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                                 (mm_interconnect_2_sysid_qsys_0_control_slave_readdata)        //                                                              .readdata
	);

	mysystem_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	mysystem_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (sys_clk_reset_source_reset),     // reset_in0.reset
		.clk            (pll_0_outclk0_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (sys_clk_reset_source_reset),         // reset_in0.reset
		.clk            (sys_clk_sys_clk_clk),                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (sys_clk_sys_clk_clk),                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
